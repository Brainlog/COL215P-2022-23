library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package data is
  type control_state is (S0, -- start state
                         S1,
                         S2,
                         S3,
                         S4,
                         S5,
                         S6,
                         S7,
                         S8,
                         S9,
                         S10,
                         S11,
                         S12,
                         S13);
end package;
